�� sr RelationInfo.��LH� I 
nbColonnesI 
nbcolonnesL 
headerPaget LPageId;L listet Ljava/util/ArrayList;L nomRelationt Ljava/lang/String;xp       sr PageId!4���]� I fileIdxI pageIdxL pageInFramet Ljava/lang/Boolean;xp        sr java.lang.Boolean� r�՜�� Z valuexpsr java.util.ArrayListx����a� I sizexp   w   sr ColInfoWS0 ���i L nomq ~ L typeq ~ xpt (Nomt VARCHAR(15)sq ~ t Prenomt VARCHAR(15)sq ~ t Aget INTEGERxt Etudiant